-------------------------------------------------------------------------------- 
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /   Vendor: Xilinx 
-- \   \   \/    Author: John F. Snow
--  \   \        Filename: $RCSfile: LCDAUX3.VHD,rcs $
--  /   /        Date Last Modified:  $Date: 2010-03-08 13:57:07-07 $
-- /___/   /\    Date Created: March 8, 2010
-- \   \  /  \ 
--  \___\/\___\ 
-- 
--
-- Revision History: 
-- $Log: LCDAUX3.VHD,rcs $
-- Revision 1.0  2010-03-08 13:57:07-07  jsnow
-- Initial release.
--
-------------------------------------------------------------------------------- 
--   
-- (c) Copyright 2010 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of,
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 
--
-------------------------------------------------------------------------------- 
--
-- Module Description:
--
-- This is the second bank of the PicoBlaze instruction ROM for the LCD control
-- module.
--------------------------------------------------------------------------------
--
-- Definition of a single port ROM for KCPSM3 program defined by lcdaux3.psm
--
-- Generated by KCPSM3 Assembler {timestamp}. 
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity lcdaux3 is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end lcdaux3;
--
architecture low_level_definition of lcdaux3 is
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  generic map ( INIT_00 => X"00090314A000540AC20100040219A0005405C10100000128A0005401C0010007",
                INIT_01 => X"C408A4F01450A0000013C440A4F8A000C440E4010000C440E401A000540FC301",
                INIT_02 => X"C440C40CA4F01450A000C44004F0000400190406040604060407145000000019",
                INIT_03 => X"E401C440040EA000C44004F000040013C4400406040604070407145000000013",
                INIT_04 => X"000E000E000EA5F0C440E40140050000C440E4010000C440E40145050000C440",
                INIT_05 => X"001904200004001900090019000E00190430000EA0000004C4400404D500000E",
                INIT_06 => X"C580A50F50722510A00000090009001D0501001D050C001D0506001D05280004",
                INIT_07 => X"A0000080A50F15F00080050E050E050E050E15F0A000001DC5C0A50FA000001D",
                INIT_08 => X"400451684003512E400250EE400150AA4000A000002C8531408585305C84450A",
                INIT_09 => X"400D5230400C5223400B520E400A5207400951FE400851C2400751AF4006518A",
                INIT_0A => X"054D002C0546006C05100067A000526340125258401152434010523F400E523B",
                INIT_0B => X"056D002C0520002C0541002C0547002C0550002C0546002C0520002C0543002C",
                INIT_0C => X"0572006C0520002C0565002C0562002C0520002C0574002C0573002C0575002C",
                INIT_0D => X"0520002C0572002C056F002C052000764F81002C0520002C0576002C0565002C",
                INIT_0E => X"05100067A000002C0572002C0565002C0568002C0567002C0569002C0568002C",
                INIT_0F => X"0520002C0574002C056E002C0565002C0572002C0572002C0575002C0543006C",
                INIT_10 => X"0541002C0547002C0550002C0546002C0520002C0543002C054D002C0546002C",
                INIT_11 => X"056F002C0569002C0573002C0569002C0576002C0565002C0572006C0520002C",
                INIT_12 => X"05100067A00000764F80002C0520002C0573002C0569002C0520002C056E002C",
                INIT_13 => X"0575002C0520002C0565002C0573002C0561002C0565002C056C002C0550006C",
                INIT_14 => X"0568002C0574006C0520002C0565002C0574002C0561002C0564002C0570002C",
                INIT_15 => X"0550002C0546002C0520002C0543002C054D002C0546002C0520002C0565002C",
                INIT_16 => X"0543002C054D002C0546006C05100067A000002C052E002C0541002C0547002C",
                INIT_17 => X"0565002C0552002C0520002C0541002C0547002C0550002C0546002C0520002C",
                INIT_18 => X"056C002C0543006C05100067A00000764F80002C0520002C053A002C0576002C",
                INIT_19 => X"0565002C056C002C0575002C0564002C056F002C056D002C0520002C056B002C",
                INIT_1A => X"0067A000026A006C0520002C0573002C0569002C0520002C15C0002C0520002C",
                INIT_1B => X"0521002C0572002C056F002C0572002C0572002C0565006C052001E5006C0510",
                INIT_1C => X"002C0575002C056D006C0520002C15F0002C052001E5006C05100067A000002C",
                INIT_1D => X"002C0579002C0574002C0520002C0565002C0562002C0520002C0574002C0573",
                INIT_1E => X"0520002C056B002C0563002C056F002C056C002C0543A000002C0565002C0570",
                INIT_1F => X"002C054EA000002C0565002C056C002C0575002C0564002C056F002C056D002C",
                INIT_20 => X"002C054EA000002C054C002C0541002C0550A000002C0543002C0553002C0554",
                INIT_21 => X"002C0565002C056B002C0563002C056F002C054C002C0520002C0574002C056F",
                INIT_22 => X"A000002C0549002C0544002C0553002C052D002C0544002C0553A000002C0564",
                INIT_23 => X"0233A000002C05410233A000002C05200227002C0547002C05334225002C0548",
                INIT_24 => X"056E002C0565002C0572002C0565002C0566002C0565002C0552A000002C0542",
                INIT_25 => X"002C0561002C0563002C056F002C054CA000002C0520002C0565002C0563002C",
                INIT_26 => X"0554528E4F00567F4D01AD03A000002C0574002C0578002C0545A000002C056C",
                INIT_27 => X"0555A00000761FE00076002C0520002C053A002C0565002C0570002C0579002C",
                INIT_28 => X"566F4E01A000002C056E002C0577002C056F002C056E002C056B002C056E002C",
                INIT_29 => X"0520A000002C0531002C054D002C0543002C054C002C0553002C0554002C0543",
                INIT_2A => X"52CB4E6052C84E5052C64E4052C14E3052C44E2052C14E1052BF4E00AEF0006C",
                INIT_2B => X"030342DB52D94ED052D74EC052D44EB052D24EA052CF4E9052DE4E8052CD4E70",
                INIT_2C => X"02E942E602E942E002FDA000032C02FD42E302FD42E602FFA000034102FF42E6",
                INIT_2D => X"42E0030EA000034102FD42E602FD42E002E9A000032C02E942E302E9A0000341",
                INIT_2E => X"0570002C0530002C0532002C0537435157462D01433C57312D01432757162D01",
                INIT_2F => X"02F442EF02F4A000002C0530002C0538002C0530002C0531A000002C0520002C",
                INIT_30 => X"057002F442F1002C0569002C0535002C0533002C0530002C053142F1002C0569",
                INIT_31 => X"002C0538002C0539002C052E002C0533002C053242F1002C0546002C0553002C",
                INIT_32 => X"002C0535002C05324320002C0534002C0532A000002C057A002C0548002C0520",
                INIT_33 => X"002C0530002C05334320002C0537002C0539002C052E002C0539002C05324320",
                INIT_34 => X"002C0534002C0539002C052E002C0539002C05354320002C0530002C05354320",
                INIT_35 => X"00000000000000000000000000000000000000004320002C0530002C05364320",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"C08000561000C081A0001000C08000671000C081A0001000C080006C1000C081",
                INIT_3E => X"1000C081A0001000C08000871000C081A0001000C080002C1000C081A0001000",
                INIT_3F => X"000000000000000000000000A0001000C080029F1000C081A0001000C080026A",    
               INITP_00 => X"B0EA8B0B0DBF3333CFFF3B82A8838E0E228FAA8F80A3EA8F02E28E2DCB72DCB4",
               INITP_01 => X"333333333B333333333333333333333333333333333B77777777777777776DDD",
               INITP_02 => X"333333333333B3333333333333333333333333333B3333333333333333333333",
               INITP_03 => X"CB333333333332CCCCCCCCCCCCCCCF3B3333333CEF33333333333333333B3333",
               INITP_04 => X"2CF33333374B332CCCCCB3333333332CECECF33CB333332CCCCCCCCCCB332CCC",
               INITP_05 => X"FECCCCB33333DF7DFBFFEFFBFFEFFFBFFDDDDDDDDDDDDDD32CCCCCCCDB333333",
               INITP_06 => X"000000000000000000000F33CCCCCF33CCF33333CCF32CCCCCCCCF333F33333C",
               INITP_07 => X"0008B28B28B28B28B28B28B20000000000000000000000000000000000000000")
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE lcdaux3.vhd
--
------------------------------------------------------------------------------------
