-------------------------------------------------------------------------------- 
--   ____  ____ 
--  /   /\/   / 
-- /___/  \  /   Vendor: Xilinx 
-- \   \   \/    Author: John F. Snow
--  \   \        Filename: $RCSfile: LCDCTRL3.VHD,rcs $
--  /   /        Date Last Modified:  $Date: 2010-03-08 13:56:05-07 $
-- /___/   /\    Date Created: March 8, 2010
-- \   \  /  \ 
--  \___\/\___\ 
-- 
--
-- Revision History: 
-- $Log: LCDCTRL3.VHD,rcs $
-- Revision 1.0  2010-03-08 13:56:05-07  jsnow
-- Initial release.
--
-------------------------------------------------------------------------------- 
--   
-- (c) Copyright 2010 Xilinx, Inc. All rights reserved.
-- 
-- This file contains confidential and proprietary information
-- of Xilinx, Inc. and is protected under U.S. and
-- international copyright and other intellectual property
-- laws.
-- 
-- DISCLAIMER
-- This disclaimer is not a license and does not grant any
-- rights to the materials distributed herewith. Except as
-- otherwise provided in a valid license issued to you by
-- Xilinx, and to the maximum extent permitted by applicable
-- law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
-- WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
-- AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
-- BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
-- INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
-- (2) Xilinx shall not be liable (whether in contract or tort,
-- including negligence, or under any other theory of,
-- liability) for any loss or damage of any kind or nature
-- related to, arising under or in connection with these
-- materials, including for any direct, or any indirect,
-- special, incidental, or consequential loss or damage
-- (including loss of data, profits, goodwill, or any type of
-- loss or damage suffered as a result of any action brought
-- by a third party) even if such damage or loss was
-- reasonably foreseeable or Xilinx had been advised of the
-- possibility of the same.
-- 
-- CRITICAL APPLICATIONS
-- Xilinx products are not designed or intended to be fail-
-- safe, or for use in any application requiring fail-safe
-- performance, such as life-support or safety devices or
-- systems, Class III medical devices, nuclear facilities,
-- applications related to the deployment of airbags, or any
-- other applications that could lead to death, personal
-- injury, or severe property or environmental damage
-- (individually and collectively, "Critical
-- Applications"). Customer assumes the sole risk and
-- liability of any use of Xilinx products in Critical
-- Applications, subject only to applicable laws and
-- regulations governing limitations on product liability.
-- 
-- THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
-- PART OF THIS FILE AT ALL TIMES. 
--
-------------------------------------------------------------------------------- 
--
-- Module Description:
--
-- This is the PicoBlaze instruction ROM for the LCD control module.
--
--------------------------------------------------------------------------------
--
-- Definition of a single port ROM for KCPSM3 program defined by lcdctrl3.psm
--
-- Generated by KCPSM3 Assembler {timestamp}. 
--
-- Standard IEEE libraries
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
--
-- The Unisim Library is used to define Xilinx primitives. It is also used during
-- simulation. The source can be viewed at %XILINX%\vhdl\src\unisims\unisim_VCOMP.vhd
--  
library unisim;
use unisim.vcomponents.all;
--
--
entity lcdctrl3 is
    Port (      address : in std_logic_vector(9 downto 0);
            instruction : out std_logic_vector(17 downto 0);
                    clk : in std_logic);
    end lcdctrl3;
--
architecture low_level_definition of lcdctrl3 is
--
begin
--
  --Instantiate the Xilinx primitive for a block RAM
  ram_1024_x_18: RAMB16_S18
  generic map ( INIT_00 => X"552A2F04551D2F02544D2F014F0000190A20016B01480137018E018E002703DC",
                INIT_01 => X"2A0414542A0214502A0114272A2040085415AF1F4F00500854392F10542F2F08",
                INIT_02 => X"2A20A00000438710052000430740051003D6A000019814802A10145C2A081458",
                INIT_03 => X"5441B0A0C03040280A205C3C0A0E402F5441B0A0C03040280A0640340A015033",
                INIT_04 => X"401503E80003A00054454610860103E2550090601070060003D0401500194039",
                INIT_05 => X"01A64D274E230F03405F4D264E220F02405F4D254E210F01405F4D244E200F00",
                INIT_06 => X"A00003F403E8000DA00003F403E8000E506C2E0850702E0454742E0251B42E01",
                INIT_07 => X"A00003E80008A00003E80009507D2E4003D0052003E8000BA00003F403E8000C",
                INIT_08 => X"052003E80012A00003E80011508D2F9003E8001003D0051003D6B0002F404F29",
                INIT_09 => X"50B24D0150AEAD071DF0548A4C62548A4D0450D14D0250C84D014C2B4D2A03D0",
                INIT_0A => X"0E600D01A00003F40D000ED050C44D0650C14D0550BD4D0450B94D0350B64D02",
                INIT_0B => X"03F40E400D00A00003F40E400D01A00003F40E50A00003F40E600D00A00003F4",
                INIT_0C => X"511A4C36511A4C3551174C0451174C03A00003F40ED00D01A00003F40EE0A000",
                INIT_0D => X"50F54D0350F24D0250EE4D0150EAAD071DF0548A4CEB51044C3051044C2F408A",
                INIT_0E => X"0EC00D00A00003F40EC00D01A00003F40E700D0051004D0650FD4D0550F94D04",
                INIT_0F => X"A00003F40E90A00003F40EA00D00A00003F40EA00D01A00003F40EB0A00003F4",
                INIT_10 => X"A00003E80E200D00548A4D0451134D0351104D02AD071DF0A00003F40E700D01",
                INIT_11 => X"55234E004E85A00003E80009A00003E80008A00003F40E200D01A00003F40E30",
                INIT_12 => X"50154F004F8A55304E004E8B401503E800040C4C4D864E834F8250154F004F84",
                INIT_13 => X"0001018E018E03E80000BC005FE04E814F80401503E800040C484D8C4E894F88",
                INIT_14 => X"4B0055514C004B854C844D864E834F824137018E018E03E80002018E018E03E8",
                INIT_15 => X"018E03E800070F4C018E018E03E80006B0005BE055585CF055584D01AD03B000",
                INIT_16 => X"4B8B4C8A4D8C4E894F884148018E018E03EE0D014E854F8403D0051003D6018E",
                INIT_17 => X"0F48018E018E03E80006B0005BE0557B5CF0557B4D01AD03B0004B0055744C00",
                INIT_18 => X"01000200416B018E018E03EE0D014E8B4F8A03D0051003D6018E018E03E80007",
                INIT_19 => X"8001B400523043000000010002004F00A000558F820155908101559180010000",
                INIT_1A => X"8531A50315F003E2055803E2055203D0051003D6A000559A8201559B8101559C",
                INIT_1B => X"000003E8000E03E8000D03E8000C03E8000BA00003E8000AA00003E2052003E2",
                INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
                INIT_3D => X"C08010001000C081A0001000C08010001000C081A0001000C08010001000C081",
                INIT_3E => X"1000C081A0001000C08010001000C081A0001000C08010001000C081A0001000",
                INIT_3F => X"000000000000000000000000A0001000C08010001000C081A0001000C0801000",    
               INITP_00 => X"B2CDCCBCBCBCDDDDC0C0C0C0F2D710FFC03BC0B36D30EF777777C3DDDDD33FFF",
               INITP_01 => X"B2C2C2CB0B0B0DDDDDDC3777DDDDB0B2C2C2CB0B0B0DDDDDDC37774332CDCCE4",
               INITP_02 => X"3F27749D003FC0CFF0FC9DD27400FF3F3F243C00D34F0034D2CB2C2CB0DDD0B0",
               INITP_03 => X"0000000000000000000000000000000033332CB343333B776400B7740FF033FC",
               INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
               INITP_07 => X"0008828828828828828828820000000000000000000000000000000000000000")
  port map(    DI => "0000000000000000",
              DIP => "00",
               EN => '1',
               WE => '0',
              SSR => '0',
              CLK => clk,
             ADDR => address,
               DO => instruction(15 downto 0),
              DOP => instruction(17 downto 16)); 
--
end low_level_definition;
--
------------------------------------------------------------------------------------
--
-- END OF FILE lcdctrl3.vhd
--
------------------------------------------------------------------------------------
